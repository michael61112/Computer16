`define not6 1
module Not6(input[5:0] in, output[5:0] out);
    assign out = ~in;
endmodule